`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:48:47 04/21/2019 
// Design Name: 
// Module Name:    vga_controller_640_60 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga_controller_640_60 (rst,pixel_clk,HS,VS,hcounter,vcounter,blank);

input rst,pixel_clk;
output HS,VS,blank;
output [10:0] hcounter,vcounter;

parameter HMAX = 800; // maxium value for the horizontal pixel counter
parameter VMAX = 525; // maxium value for the vertical pixel counter
parameter HLINES = 640; // total number of visible columns
parameter HFP = 648; // value for the horizontal counter where front porch ends
parameter HSP = 744; // value for the horizontal counter where the synch pulse ends
parameter VLINES = 480; // total number of visible lines
parameter VFP = 482; // value for the vertical counter where the frone proch ends
parameter VSP = 484; // value for the vertical counter where the synch pulse ends
parameter SPP = 0;


wire video_enable;
reg HS,VS,blank;
reg [10:0] hcounter,vcounter;

always@(posedge pixel_clk)begin
blank <= ~video_enable; end

always@(posedge pixel_clk)begin
    if(rst == 1)
	   hcounter <= 0;
    else if (hcounter == HMAX)
	   hcounter <= 0;
    else
	   hcounter <= hcounter + 1;
end

always@(posedge pixel_clk)begin
    if(rst == 1)
	   vcounter <=0;
    else if(hcounter == HMAX) begin
      if(vcounter == VMAX)
		  vcounter <= 0;
      else
		  vcounter <= vcounter + 1;
		end
end

always@(posedge pixel_clk)begin
if(hcounter >=HFP && hcounter < HSP) HS <= SPP;
else HS <= ~SPP; end

always@(posedge pixel_clk)begin
if(vcounter >=VFP && vcounter <VSP) VS <= SPP;
else VS <= ~SPP; end

assign video_enable = (hcounter < HLINES && vcounter < VLINES)? 1'b1:1'b0;

endmodule
